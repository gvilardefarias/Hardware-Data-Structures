`define CLK_PERIOD 10
